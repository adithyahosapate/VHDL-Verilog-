

module fulladder (sum,c1,a,b,c);

output sum,c1;
input a,b,c;




assign sum=()
assign c1=(b&&c);

endmodule






